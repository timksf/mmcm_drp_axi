package GLBL;

import "BVI" glbl = 
module vMkGLBL(Empty);
    default_clock no_clock;
    default_reset no_reset;
endmodule

endpackage